library verilog;
use verilog.vl_types.all;
entity APB_Protocol_tb is
end APB_Protocol_tb;
